CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 457 276
42991634 0
0
6 Title:
5 Name:
0
0
0
42
13 Logic Switch~
5 44 191 0 1 11
0 16
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9993 0 0
2
38782 0
0
13 Logic Switch~
5 45 157 0 1 11
0 4
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
446 0 0
2
38782 1
0
13 Logic Switch~
5 46 126 0 1 11
0 15
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9386 0 0
2
38782 2
0
13 Logic Switch~
5 46 100 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
349 0 0
2
38782 3
0
9 CC 7-Seg~
183 1538 293 0 17 19
10 11 7 8 10 9 6 5 43 2
1 1 1 1 1 1 0 2
0
0 0 21360 0
5 REDCC
16 -41 51 -33
5 DISP2
14 -52 49 -44
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4860 0 0
2
38782 4
0
8 2-In OR~
219 157 337 0 3 22
0 13 12 11
0
0 0 352 0
6 74LS32
-21 -24 21 -16
4 U11C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
3914 0 0
2
38782 5
0
8 2-In OR~
219 94 346 0 3 22
0 14 4 12
0
0 0 2400 0
6 74LS32
-21 -24 21 -16
4 U11B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
3367 0 0
2
38782 6
0
6 74266~
219 99 300 0 3 22
0 16 15 13
0
0 0 2400 0
7 74LS266
-24 -24 25 -16
4 U12B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
4507 0 0
2
38782 7
0
9 Inverter~
13 214 314 0 2 22
0 15 17
0
0 0 2400 270
6 74LS04
-16 -43 26 -35
3 U9B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
6934 0 0
2
38782 8
0
6 74266~
219 291 300 0 3 22
0 16 4 18
0
0 0 2400 0
7 74LS266
-24 -24 25 -16
4 U12A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
6670 0 0
2
38782 9
0
8 2-In OR~
219 293 354 0 3 22
0 17 14 19
0
0 0 2400 0
6 74LS32
-21 -24 21 -16
4 U11A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3474 0 0
2
38782 10
0
8 2-In OR~
219 347 326 0 3 22
0 18 19 7
0
0 0 2400 0
6 74LS32
-21 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
733 0 0
2
38782 11
0
8 4-In OR~
219 526 341 0 5 22
0 16 3 15 14 8
0
0 0 2400 0
4 4072
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
3698 0 0
2
38782 12
0
9 Inverter~
13 426 311 0 2 22
0 4 3
0
0 0 2400 270
6 74LS04
-21 -19 21 -11
3 U9A
20 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
3625 0 0
2
38782 13
0
9 2-In AND~
219 1168 299 0 3 22
0 15 21 20
0
0 0 2400 0
6 74LS08
-21 -24 21 -16
3 U7C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3909 0 0
2
38782 14
0
8 3-In OR~
219 1225 332 0 4 22
0 20 22 14 6
0
0 0 2400 0
4 4075
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 8 0
1 U
8542 0 0
2
38782 15
0
8 2-In OR~
219 1111 391 0 3 22
0 21 15 23
0
0 0 2400 0
6 74LS32
-21 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
8460 0 0
2
38782 16
0
9 2-In AND~
219 1178 343 0 3 22
0 24 23 22
0
0 0 2400 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3790 0 0
2
38782 17
0
9 Inverter~
13 1110 263 0 2 22
0 4 24
0
0 0 2400 270
6 74LS04
-21 -19 21 -11
3 U6F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 6 0
1 U
435 0 0
2
38782 18
0
9 Inverter~
13 1311 316 0 2 22
0 14 25
0
0 0 2144 270
6 74LS04
-21 -19 21 -11
3 U6E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 6 0
1 U
7502 0 0
2
38782 19
0
8 4-In OR~
219 1464 336 0 5 22
0 14 27 28 26 5
0
0 0 2400 0
4 4072
-14 -24 14 -16
3 U3B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
4348 0 0
2
38782 20
0
9 Inverter~
13 1296 295 0 2 22
0 16 29
0
0 0 2144 270
6 74LS04
-21 -19 21 -11
3 U6D
20 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
3505 0 0
2
38782 21
0
9 Inverter~
13 1325 294 0 2 22
0 4 30
0
0 0 2144 270
6 74LS04
-21 -19 21 -11
3 U6C
20 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
820 0 0
2
38782 22
0
5 7415~
219 1393 350 0 4 22
0 4 31 25 26
0
0 0 2400 0
6 74LS15
-21 -28 21 -20
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 5 0
1 U
8602 0 0
2
38782 23
0
9 2-In AND~
219 1388 406 0 3 22
0 29 4 27
0
0 0 2400 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3609 0 0
2
38782 24
0
9 2-In AND~
219 1395 302 0 3 22
0 15 30 28
0
0 0 2400 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3752 0 0
2
38782 25
0
9 Inverter~
13 1341 327 0 2 22
0 15 31
0
0 0 2144 270
6 74LS04
-21 -19 21 -11
3 U6B
20 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
8387 0 0
2
38782 26
0
9 Inverter~
13 1068 263 0 2 22
0 16 21
0
0 0 2400 270
6 74LS04
-21 -19 21 -11
3 U6A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
4723 0 0
2
38782 27
0
9 2-In AND~
219 1036 362 0 3 22
0 32 33 9
0
0 0 2400 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5406 0 0
2
38782 28
0
9 Inverter~
13 975 267 0 2 22
0 15 34
0
0 0 2400 270
6 74LS04
-21 -19 21 -11
3 U2F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
5782 0 0
2
38782 29
0
9 Inverter~
13 925 267 0 2 22
0 16 32
0
0 0 2400 270
6 74LS04
-21 -19 21 -11
3 U2E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
8264 0 0
2
38782 30
0
8 2-In OR~
219 994 324 0 3 22
0 4 34 33
0
0 0 2400 0
6 74LS32
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3817 0 0
2
38782 31
0
9 2-In AND~
219 786 358 0 3 22
0 36 4 35
0
0 0 2400 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3315 0 0
2
38782 32
0
9 Inverter~
13 700 406 0 2 22
0 4 37
0
0 0 2400 0
6 74LS04
-21 -19 21 -11
3 U2D
20 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
3438 0 0
2
38782 33
0
5 7415~
219 776 397 0 4 22
0 15 16 37 38
0
0 0 2400 0
6 74LS15
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 5 0
1 U
9921 0 0
2
38782 34
0
9 Inverter~
13 721 322 0 2 22
0 15 39
0
0 0 2400 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
9469 0 0
2
38782 35
0
9 Inverter~
13 723 457 0 2 22
0 15 40
0
0 0 2400 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3716 0 0
2
38782 36
0
9 2-In AND~
219 787 448 0 3 22
0 42 40 41
0
0 0 2400 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3768 0 0
2
38782 37
0
8 4-In OR~
219 868 362 0 5 22
0 38 35 41 14 10
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
3830 0 0
2
38782 38
0
9 Inverter~
13 718 301 0 2 22
0 16 42
0
0 0 2400 0
6 74LS04
-21 -19 21 -11
3 U2A
20 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3377 0 0
2
38782 39
0
8 2-In OR~
219 779 310 0 3 22
0 42 39 36
0
0 0 2400 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3102 0 0
2
38782 40
0
7 Ground~
168 1590 349 0 1 3
0 2
0
0 0 55904 0
0
4 GND1
4 -11 32 -3
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7960 0 0
2
38782 41
0
75
2 2 3 0 0 8320 0 14 13 0 0 3
429 329
429 337
509 337
0 1 4 0 0 8192 0 0 24 47 0 3
1277 339
1277 341
1369 341
5 7 5 0 0 12432 0 21 5 0 0 4
1497 336
1497 419
1553 419
1553 329
4 6 6 0 0 8320 0 16 5 0 0 4
1258 332
1258 432
1547 432
1547 329
2 0 4 0 0 4096 0 33 0 0 72 2
762 367
647 367
2 3 7 0 0 8320 0 5 12 0 0 5
1523 329
1523 467
393 467
393 326
380 326
5 3 8 0 0 8320 0 13 5 0 0 4
559 341
559 507
1529 507
1529 329
3 5 9 0 0 8320 0 29 5 0 0 4
1057 362
1057 451
1541 451
1541 329
5 4 10 0 0 8320 0 39 5 0 0 4
901 362
901 488
1535 488
1535 329
9 1 2 0 0 12416 0 5 42 0 0 4
1538 251
1538 218
1590 218
1590 343
3 1 11 0 0 8320 0 6 5 0 0 4
190 337
190 478
1517 478
1517 329
3 2 12 0 0 4224 0 7 6 0 0 2
127 346
144 346
3 1 13 0 0 4224 0 8 6 0 0 3
138 300
138 328
144 328
1 1 14 0 0 8192 0 4 7 0 0 4
58 100
63 100
63 337
81 337
0 2 4 0 0 4096 0 0 7 71 0 3
72 157
72 355
81 355
0 2 15 0 0 4096 0 0 8 75 0 3
66 126
66 309
83 309
0 1 16 0 0 4096 0 0 8 69 0 3
77 191
77 291
83 291
2 1 17 0 0 8320 0 9 11 0 0 3
217 332
217 345
280 345
0 1 15 0 0 0 0 0 9 75 0 2
217 126
217 296
3 1 18 0 0 4224 0 10 12 0 0 3
330 300
330 317
334 317
0 2 4 0 0 0 0 0 10 71 0 3
233 157
233 309
275 309
0 1 16 0 0 0 0 0 10 69 0 3
254 191
254 291
275 291
3 2 19 0 0 8320 0 11 12 0 0 4
326 354
330 354
330 335
334 335
0 2 14 0 0 4096 0 0 11 70 0 3
198 100
198 363
280 363
0 4 14 0 0 0 0 0 13 70 0 3
399 100
399 355
509 355
0 3 15 0 0 4096 0 0 13 75 0 3
413 126
413 346
509 346
0 1 16 0 0 4096 0 0 13 69 0 3
471 191
471 328
509 328
0 1 4 0 0 0 0 0 14 71 0 2
429 157
429 293
3 1 20 0 0 8320 0 15 16 0 0 4
1189 299
1204 299
1204 323
1212 323
0 2 21 0 0 4096 0 0 15 35 0 2
1071 308
1144 308
0 1 15 0 0 0 0 0 15 36 0 4
1090 288
1136 288
1136 290
1144 290
3 2 22 0 0 8320 0 18 16 0 0 4
1199 343
1204 343
1204 332
1213 332
0 3 14 0 0 0 0 0 16 70 0 3
1208 100
1208 341
1212 341
3 2 23 0 0 8320 0 17 18 0 0 4
1144 391
1148 391
1148 352
1154 352
1 2 21 0 0 8320 0 17 28 0 0 3
1098 382
1071 382
1071 281
0 2 15 0 0 4096 0 0 17 75 0 3
1090 126
1090 400
1098 400
2 1 24 0 0 4224 0 19 18 0 0 3
1113 281
1113 334
1154 334
0 1 4 0 0 0 0 0 19 71 0 4
1110 157
1110 237
1113 237
1113 245
2 3 25 0 0 8320 0 20 24 0 0 3
1314 334
1314 359
1369 359
4 4 26 0 0 4224 0 24 21 0 0 2
1414 350
1447 350
3 2 27 0 0 8320 0 25 21 0 0 4
1409 406
1434 406
1434 332
1447 332
3 3 28 0 0 8320 0 26 21 0 0 4
1416 302
1439 302
1439 341
1447 341
0 1 14 0 0 0 0 0 21 70 0 5
1314 100
1427 100
1427 324
1447 324
1447 323
2 1 29 0 0 8320 0 22 25 0 0 4
1299 313
1285 313
1285 397
1364 397
2 2 30 0 0 12416 0 23 26 0 0 5
1328 312
1328 370
1358 370
1358 311
1371 311
2 2 31 0 0 8320 0 27 24 0 0 3
1344 345
1344 350
1369 350
0 2 4 0 0 8192 0 0 25 71 0 4
1274 157
1277 157
1277 415
1364 415
0 1 15 0 0 0 0 0 27 75 0 2
1344 126
1344 309
0 1 16 0 0 0 0 0 28 69 0 2
1071 191
1071 245
2 1 32 0 0 8320 0 31 29 0 0 3
928 285
928 353
1012 353
3 2 33 0 0 16512 0 32 29 0 0 6
1027 324
1031 324
1031 343
1007 343
1007 371
1012 371
2 2 34 0 0 4224 0 30 32 0 0 3
978 285
978 333
981 333
0 1 15 0 0 0 0 0 30 75 0 4
977 126
977 241
978 241
978 249
0 1 16 0 0 0 0 0 31 69 0 2
928 191
928 249
0 1 4 0 0 0 0 0 32 71 0 3
951 157
951 315
981 315
3 2 35 0 0 4224 0 33 39 0 0 2
807 358
851 358
1 3 36 0 0 8320 0 33 41 0 0 6
762 349
761 349
761 290
820 290
820 310
812 310
3 2 37 0 0 4224 0 35 34 0 0 2
752 406
721 406
1 4 38 0 0 8320 0 39 35 0 0 4
851 349
805 349
805 397
797 397
0 1 15 0 0 0 0 0 35 74 0 2
635 388
752 388
0 2 16 0 0 0 0 0 35 73 0 5
661 300
661 429
739 429
739 397
752 397
2 2 39 0 0 4224 0 36 41 0 0 4
742 322
758 322
758 319
766 319
0 1 15 0 0 0 0 0 36 74 0 2
635 322
706 322
2 2 40 0 0 4224 0 37 38 0 0 2
744 457
763 457
3 3 41 0 0 8320 0 38 39 0 0 4
808 448
833 448
833 367
851 367
2 1 42 0 0 8320 0 40 38 0 0 4
739 301
745 301
745 439
763 439
0 4 14 0 0 0 0 0 39 70 0 7
614 100
614 360
755 360
755 331
843 331
843 376
851 376
2 1 42 0 0 0 0 40 41 0 0 2
739 301
766 301
1 1 16 0 0 8320 0 22 1 0 0 3
1299 277
1299 191
56 191
1 1 14 0 0 8320 0 20 4 0 0 3
1314 298
1314 100
58 100
1 1 4 0 0 8320 0 23 2 0 0 3
1328 276
1328 157
57 157
0 1 4 0 0 0 0 0 34 71 0 3
647 157
647 406
685 406
0 1 16 0 0 0 0 0 40 69 0 3
661 191
661 301
703 301
0 1 15 0 0 4096 0 0 37 75 0 3
635 126
635 457
708 457
1 1 15 0 0 4224 0 3 26 0 0 4
58 126
1363 126
1363 293
1371 293
2
-21 0 0 0 700 0 0 0 0 1 2 1 49
8 Fixedsys
0 0 0 34
510 43 826 64
514 47 821 62
34 DECODIFICADOR DE BINARIO A DECIMAL
-27 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 38
208 7 827 54
213 11 821 42
38 UNIVERSIDAD TECNOLOGICA DE EL SALVADOR
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
