CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
150 0 30 100 9
0 66 1024 740
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
72 C:\ARCHIVOS DE PROGRAMA\MICROCODE ENGINEERING\CIRCUITMAKER 6 PRO\BOM.DAT
0 7
0 66 1024 740
177209362 0
0
6 Title:
5 Name:
0
0
0
33
13 Logic Switch~
5 1082 725 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 508 986 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 492 808 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 469 778 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 326 757 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 312 717 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 305 867 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 366 51 0 1 11
0 39
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3747 0 0
0
0
5 4011~
219 1314 996 0 3 21
0 11 10 6
0
0 0 624 512
4 4011
-7 -24 21 -16
4 U11D
-11 -25 17 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 2 0
1 U
3549 0 0
0
0
5 4011~
219 1316 950 0 3 21
0 11 9 5
0
0 0 624 512
4 4011
-7 -24 21 -16
4 U11C
-11 -25 17 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 2 0
1 U
7931 0 0
0
0
5 4011~
219 1313 897 0 3 21
0 11 8 4
0
0 0 624 512
4 4011
-7 -24 21 -16
4 U11B
-11 -25 17 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 2 0
1 U
9325 0 0
0
0
5 4011~
219 1308 833 0 3 21
0 11 7 3
0
0 0 624 512
4 4011
-7 -24 21 -16
4 U11A
-11 -25 17 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -1610612604
65 0 0 0 4 1 2 0
1 U
8903 0 0
0
0
8 Hex Key~
166 1357 737 0 11 12
0 10 9 8 7 0 0 0 0 0
7 55
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
3834 0 0
0
0
2 +V
167 1141 789 0 1 3
0 12
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3363 0 0
0
0
7 Ground~
168 1007 791 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7668 0 0
0
0
8 Hex Key~
166 939 799 0 11 12
0 16 15 14 13 0 0 0 0 0
6 54
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
4718 0 0
0
0
12 Hex Display~
7 1214 806 0 18 19
10 6 5 4 3 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3874 0 0
0
0
6 1K RAM
79 1110 883 0 20 41
0 2 2 2 2 2 2 13 14 15
16 50 51 52 53 3 4 5 6 12
11
0
0 0 13040 0
5 RAM1K
-17 -19 18 -11
3 U10
-11 -70 10 -62
0
15 DVCC=22;DGND=11
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 -1610612668
65 0 0 512 0 0 0 0
1 U
6671 0 0
0
0
7 Ground~
168 275 264 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3789 0 0
0
0
7 74LS160
124 154 350 0 14 29
0 54 55 56 57 58 59 60 61 62
63 25 26 27 28
0
0 0 13040 0
8 74LS160A
-27 -51 29 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 -1610612592
65 0 0 512 1 0 0 0
1 U
4871 0 0
0
0
12 Hex Display~
7 634 825 0 16 19
10 38 37 36 35 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3750 0 0
0
0
7 74LS161
96 461 888 0 14 29
0 29 30 34 64 65 66 67 31 32
33 35 36 37 38
0
0 0 13040 0
8 74LS161A
-28 -60 28 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 -1610612592
65 0 0 512 1 0 0 0
1 U
8778 0 0
0
0
7 Ground~
168 698 231 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
538 0 0
0
0
5 7405~
219 811 180 0 2 21
0 39 40
0
0 0 624 270
6 74LS05
-21 -24 21 -16
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 -1610612604
65 0 0 0 6 1 1 0
1 U
6843 0 0
0
0
8 Hex Key~
166 639 103 0 11 12
0 24 23 22 21 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
3136 0 0
0
0
12 Hex Display~
7 1277 426 0 16 19
10 44 43 42 41 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
5950 0 0
0
0
4 4042
219 1147 195 0 14 29
0 68 69 70 71 72 73 74 75 76
77 78 79 80 81
0
0 0 13040 0
4 4042
-14 -60 14 -52
2 U7
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 14 13 7 4 6 5 3 2 9
10 12 11 15 1 14 13 7 4 6
5 3 2 9 10 12 11 15 1 -1610612592
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
7 74LS160
124 1157 522 0 14 29
0 82 83 45 84 85 86 87 88 89
90 41 42 43 44
0
0 0 13040 0
8 74LS160A
-27 -51 29 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 -1610612592
65 0 0 512 1 0 0 0
1 U
6828 0 0
0
0
6 74LS85
106 948 480 0 14 29
0 46 47 48 49 17 18 19 20 91
92 93 94 45 95
0
0 0 13296 0
6 74LS85
-21 -52 21 -44
2 U5
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 -1610612676
65 0 0 512 1 0 0 0
1 U
6735 0 0
0
0
7 Ground~
168 620 382 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8365 0 0
0
0
7 74LS245
64 721 431 0 18 37
0 96 97 98 99 21 22 23 24 100
101 102 17 103 18 19 20 2 39
0
0 0 13040 0
7 74LS245
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
4132 0 0
0
0
7 74LS245
64 743 298 0 18 37
0 104 105 106 107 21 22 23 24 108
109 110 111 46 47 48 49 2 40
0
0 0 13040 0
7 74LS245
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
4551 0 0
0
0
6 1K RAM
79 322 341 0 20 41
0 2 2 2 2 2 2 25 26 27
28 112 113 114 115 17 18 19 20 116
39
0
0 0 13040 0
5 RAM1K
-17 -19 18 -11
2 U4
-7 -70 7 -62
0
15 DVCC=22;DGND=11
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 -1610612676
65 0 0 512 0 0 0 0
1 U
3635 0 0
0
0
79
3 0 3 0 0 4096 0 12 0 0 25 4
1283 833
1235 833
1235 853
1205 853
3 0 4 0 0 4224 0 11 0 0 26 3
1288 897
1174 897
1174 910
3 0 5 0 0 4224 0 10 0 0 27 3
1291 950
1169 950
1169 919
3 0 6 0 0 4224 0 9 0 0 28 3
1289 996
1162 996
1162 928
4 2 7 0 0 4224 0 13 12 0 0 3
1348 761
1348 842
1334 842
3 2 8 0 0 4224 0 13 11 0 0 3
1354 761
1354 906
1339 906
2 2 9 0 0 4224 0 13 10 0 0 3
1360 761
1360 959
1342 959
1 2 10 0 0 4224 0 13 9 0 0 3
1366 761
1366 1005
1340 1005
0 1 11 0 0 8192 0 0 9 10 0 4
1351 940
1349 940
1349 987
1340 987
0 1 11 0 0 0 0 0 10 11 0 4
1348 896
1351 896
1351 941
1342 941
0 1 11 0 0 8192 0 0 11 12 0 6
1340 819
1280 819
1280 917
1348 917
1348 888
1339 888
0 1 11 0 0 4224 0 0 12 14 0 6
1156 735
1337 735
1337 814
1340 814
1340 824
1334 824
1 19 12 0 0 12416 0 14 18 0 0 5
1141 798
1141 819
1142 819
1142 847
1148 847
1 20 11 0 0 128 0 1 18 0 0 4
1094 725
1156 725
1156 856
1148 856
1 0 2 0 0 8192 0 18 0 0 20 3
1078 847
1078 848
1070 848
2 0 2 0 0 0 0 18 0 0 20 3
1078 856
1078 857
1070 857
3 0 2 0 0 0 0 18 0 0 20 3
1078 865
1078 867
1070 867
4 0 2 0 0 0 0 18 0 0 20 3
1078 874
1078 875
1070 875
5 0 2 0 0 0 0 18 0 0 20 3
1078 883
1078 884
1070 884
1 6 2 0 0 12416 0 15 18 0 0 5
1007 785
1007 781
1070 781
1070 892
1078 892
4 7 13 0 0 8320 0 16 18 0 0 3
930 823
930 901
1078 901
3 8 14 0 0 8320 0 16 18 0 0 3
936 823
936 910
1078 910
2 9 15 0 0 8320 0 16 18 0 0 3
942 823
942 919
1078 919
1 10 16 0 0 8320 0 16 18 0 0 3
948 823
948 928
1078 928
4 15 3 0 0 4224 0 17 18 0 0 3
1205 830
1205 901
1142 901
3 16 4 0 0 128 0 17 18 0 0 3
1211 830
1211 910
1142 910
2 17 5 0 0 128 0 17 18 0 0 3
1217 830
1217 919
1142 919
1 18 6 0 0 128 0 17 18 0 0 3
1223 830
1223 928
1142 928
1 0 2 0 0 0 0 33 0 0 34 2
290 305
282 305
2 0 2 0 0 0 0 33 0 0 34 2
290 314
282 314
3 0 2 0 0 0 0 33 0 0 34 3
290 323
290 325
282 325
4 0 2 0 0 0 0 33 0 0 34 3
290 332
290 333
282 333
5 0 2 0 0 0 0 33 0 0 34 2
290 341
282 341
1 6 2 0 0 0 0 19 33 0 0 7
275 258
275 254
289 254
289 277
282 277
282 350
290 350
12 0 17 0 0 8192 0 31 0 0 43 3
753 431
780 431
780 494
14 0 18 0 0 8192 0 31 0 0 44 3
753 449
773 449
773 500
15 0 19 0 0 8192 0 31 0 0 45 3
753 458
766 458
766 507
16 0 20 0 0 8192 0 31 0 0 46 3
753 467
757 467
757 516
5 0 21 0 0 8192 0 31 0 0 66 3
689 440
655 440
655 307
6 0 22 0 0 8192 0 31 0 0 67 3
689 449
662 449
662 316
7 0 23 0 0 8192 0 31 0 0 68 3
689 458
671 458
671 325
8 0 24 0 0 8192 0 31 0 0 69 3
689 467
679 467
679 334
15 5 17 0 0 8320 0 33 29 0 0 5
354 359
354 494
908 494
908 489
916 489
16 6 18 0 0 8320 0 33 29 0 0 5
354 368
354 500
908 500
908 498
916 498
17 7 19 0 0 8320 0 33 29 0 0 3
354 377
354 507
916 507
18 8 20 0 0 16512 0 33 29 0 0 5
354 386
354 517
607 517
607 516
916 516
11 7 25 0 0 4224 0 20 33 0 0 2
186 359
290 359
12 8 26 0 0 4224 0 20 33 0 0 2
186 368
290 368
13 9 27 0 0 4224 0 20 33 0 0 2
186 377
290 377
14 10 28 0 0 4224 0 20 33 0 0 2
186 386
290 386
1 1 29 0 0 8320 0 6 22 0 0 4
324 717
421 717
421 852
429 852
1 2 30 0 0 8320 0 5 22 0 0 4
338 757
421 757
421 861
429 861
1 8 31 0 0 8320 0 4 22 0 0 4
481 778
510 778
510 852
499 852
1 9 32 0 0 8320 0 3 22 0 0 4
504 808
509 808
509 861
499 861
1 10 33 0 0 8320 0 2 22 0 0 4
520 986
525 986
525 888
493 888
1 3 34 0 0 4224 0 7 22 0 0 4
317 867
421 867
421 870
429 870
4 11 35 0 0 8320 0 21 22 0 0 3
625 849
625 897
493 897
3 12 36 0 0 8320 0 21 22 0 0 3
631 849
631 906
493 906
2 13 37 0 0 8320 0 21 22 0 0 3
637 849
637 915
493 915
1 14 38 0 0 8320 0 21 22 0 0 3
643 849
643 924
493 924
1 17 2 0 0 128 0 23 32 0 0 5
698 225
698 221
697 221
697 262
705 262
0 20 39 0 0 4096 0 0 33 65 0 3
412 51
412 314
360 314
0 18 39 0 0 0 0 0 31 65 0 4
814 140
854 140
854 395
753 395
2 18 40 0 0 4224 0 24 32 0 0 3
814 198
814 262
775 262
1 1 39 0 0 4224 0 8 24 0 0 3
378 51
814 51
814 162
4 5 21 0 0 4224 0 25 32 0 0 3
630 127
630 307
711 307
3 6 22 0 0 4224 0 25 32 0 0 3
636 127
636 316
711 316
2 7 23 0 0 4224 0 25 32 0 0 3
642 127
642 325
711 325
1 8 24 0 0 4224 0 25 32 0 0 3
648 127
648 334
711 334
4 11 41 0 0 4224 0 26 28 0 0 3
1268 450
1268 531
1189 531
3 12 42 0 0 4224 0 26 28 0 0 3
1274 450
1274 540
1189 540
2 13 43 0 0 4224 0 26 28 0 0 3
1280 450
1280 549
1189 549
1 14 44 0 0 4224 0 26 28 0 0 3
1286 450
1286 558
1189 558
13 3 45 0 0 4224 0 29 28 0 0 4
980 507
1111 507
1111 513
1125 513
1 13 46 0 0 8320 0 29 32 0 0 4
916 453
783 453
783 307
775 307
2 14 47 0 0 8320 0 29 32 0 0 4
916 462
783 462
783 316
775 316
3 15 48 0 0 8320 0 29 32 0 0 4
916 471
783 471
783 325
775 325
4 16 49 0 0 8320 0 29 32 0 0 4
916 480
783 480
783 334
775 334
1 17 2 0 0 128 0 30 31 0 0 4
620 376
618 376
618 395
683 395
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
