CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
150 0 30 100 10
176 83 798 549
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 457 276
42991634 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 56 66 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3752 0 0
2
38793.6 0
0
13 Logic Switch~
5 55 114 0 1 11
0 39
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7343 0 0
2
38793.6 1
0
13 Logic Switch~
5 56 160 0 1 11
0 40
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7856 0 0
2
38793.6 2
0
13 Logic Switch~
5 54 208 0 1 11
0 41
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7796 0 0
2
38793.6 3
0
13 Logic Switch~
5 55 257 0 1 11
0 42
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7567 0 0
2
38793.6 4
0
13 Logic Switch~
5 53 309 0 1 11
0 43
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8638 0 0
2
38793.6 5
0
13 Logic Switch~
5 56 355 0 1 11
0 44
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
321 0 0
2
38793.6 6
0
13 Logic Switch~
5 54 402 0 1 11
0 45
0
0 0 21360 0
2 0V
-7 -16 7 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5556 0 0
2
38793.6 7
0
2 +V
167 1068 35 0 1 3
0 3
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7958 0 0
2
38793.6 8
0
9 CA 7-Seg~
184 1068 116 0 18 19
10 4 5 6 7 8 9 10 46 3
0 0 0 0 0 0 0 2 1
0
0 0 21344 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
377 0 0
2
38793.6 9
0
6 74LS47
187 949 213 0 14 29
0 14 13 12 11 47 48 10 9 8
7 6 5 4 49
0
0 0 4848 0
6 74LS47
-21 -60 21 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5955 0 0
2
38793.6 10
0
7 74LS157
122 809 211 0 14 29
0 23 22 18 21 17 20 16 19 15
2 14 13 12 11
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3291 0 0
2
38793.6 11
0
5 4049~
219 624 253 0 2 22
0 26 27
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 1 0
1 U
8824 0 0
2
38793.6 12
0
5 4081~
219 686 223 0 3 22
0 28 27 23
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
7556 0 0
2
38793.6 13
0
5 4071~
219 556 253 0 3 22
0 25 24 26
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3269 0 0
2
38793.6 14
0
7 Ground~
168 399 505 0 1 3
0 2
0
0 0 49264 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9627 0 0
2
38793.6 15
0
12 Hex Display~
7 220 48 0 18 19
10 30 31 32 33 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5470 0 0
2
38793.6 16
0
6 74LS85
106 455 224 0 14 29
0 33 32 31 30 2 29 2 29 50
51 52 28 25 24
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U5
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7104 0 0
2
38793.6 17
0
6 74LS83
105 556 356 0 14 29
0 33 32 31 30 2 2 2 29 2
18 17 16 15 53
0
0 0 4848 0
7 74LS83A
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
5265 0 0
2
38793.6 18
0
6 74LS83
105 560 76 0 14 29
0 33 32 31 30 2 2 29 2 2
22 21 20 19 54
0
0 0 4848 0
7 74LS83A
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
472 0 0
2
38793.6 19
0
5 4049~
219 289 283 0 2 22
0 34 30
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 1 0
1 U
3415 0 0
2
38793.6 20
0
5 4049~
219 289 248 0 2 22
0 35 31
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
52 0 0
2
38793.6 21
0
5 4049~
219 288 210 0 2 22
0 36 32
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
4810 0 0
2
38793.6 22
0
5 4049~
219 287 176 0 2 22
0 37 33
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
3794 0 0
2
38793.6 23
0
5 74147
219 198 225 0 13 27
0 55 38 39 40 41 42 43 44 45
34 35 36 37
0
0 0 4848 0
5 74147
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
121 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
27

0 10 5 4 3 2 1 13 12 11
9 7 6 14 10 5 4 3 2 1
13 12 11 9 7 6 14 0
65 0 0 512 1 0 0 0
1 U
4110 0 0
2
38793.6 24
0
68
9 1 3 0 0 4224 0 10 9 0 0 2
1068 80
1068 44
13 1 4 0 0 8320 0 11 10 0 0 3
987 231
1047 231
1047 152
12 2 5 0 0 8320 0 11 10 0 0 3
987 222
1053 222
1053 152
11 3 6 0 0 4224 0 11 10 0 0 3
987 213
1059 213
1059 152
10 4 7 0 0 4224 0 11 10 0 0 3
987 204
1065 204
1065 152
9 5 8 0 0 4224 0 11 10 0 0 3
987 195
1071 195
1071 152
8 6 9 0 0 4224 0 11 10 0 0 3
987 186
1077 186
1077 152
7 7 10 0 0 4224 0 11 10 0 0 3
987 177
1083 177
1083 152
4 14 11 0 0 4224 0 11 12 0 0 4
917 204
859 204
859 247
841 247
3 13 12 0 0 4224 0 11 12 0 0 4
917 195
849 195
849 229
841 229
2 12 13 0 0 4224 0 11 12 0 0 4
917 186
854 186
854 211
841 211
1 11 14 0 0 4224 0 11 12 0 0 4
917 177
849 177
849 193
841 193
10 0 2 0 0 12288 0 12 0 0 40 4
771 256
649 256
649 290
399 290
13 9 15 0 0 4224 0 19 12 0 0 4
588 374
748 374
748 247
777 247
12 7 16 0 0 4224 0 19 12 0 0 4
588 365
763 365
763 229
777 229
11 5 17 0 0 4224 0 19 12 0 0 4
588 356
753 356
753 211
777 211
10 3 18 0 0 4224 0 19 12 0 0 4
588 347
758 347
758 193
777 193
13 8 19 0 0 4224 0 20 12 0 0 4
592 94
743 94
743 238
777 238
12 6 20 0 0 4224 0 20 12 0 0 4
592 85
748 85
748 220
777 220
11 4 21 0 0 4224 0 20 12 0 0 4
592 76
753 76
753 202
777 202
10 2 22 0 0 4224 0 20 12 0 0 4
592 67
758 67
758 184
777 184
3 1 23 0 0 4224 0 14 12 0 0 4
707 223
763 223
763 175
777 175
2 14 24 0 0 4224 0 15 18 0 0 4
543 262
502 262
502 260
487 260
1 13 25 0 0 4224 0 15 18 0 0 4
543 244
500 244
500 251
487 251
1 3 26 0 0 4224 0 13 15 0 0 2
609 253
589 253
2 2 27 0 0 8320 0 14 13 0 0 4
662 232
655 232
655 253
645 253
1 12 28 0 0 12416 0 14 18 0 0 6
662 214
644 214
644 231
495 231
495 242
487 242
5 0 2 0 0 0 0 19 0 0 31 2
524 356
478 356
6 0 2 0 0 0 0 19 0 0 31 3
524 365
486 365
486 401
7 0 2 0 0 0 0 19 0 0 31 3
524 374
493 374
493 401
9 0 2 0 0 0 0 19 0 0 35 3
524 401
478 401
478 309
8 0 2 0 0 0 0 20 0 0 35 4
528 103
508 103
508 180
520 180
6 0 2 0 0 0 0 20 0 0 35 4
528 85
513 85
513 150
520 150
5 0 2 0 0 0 0 20 0 0 35 4
528 76
523 76
523 121
520 121
0 9 2 0 0 0 0 0 20 40 0 4
399 309
520 309
520 121
528 121
7 0 29 0 0 8320 0 20 0 0 37 3
528 94
419 94
419 242
6 0 29 0 0 0 0 18 0 0 38 3
423 242
419 242
419 266
8 8 29 0 0 0 0 18 19 0 0 4
423 260
419 260
419 383
524 383
7 0 2 0 0 0 0 18 0 0 40 2
423 251
399 251
5 1 2 0 0 8320 0 18 16 0 0 3
423 233
399 233
399 499
0 1 30 0 0 4096 0 0 17 49 0 3
359 80
229 80
229 72
0 2 31 0 0 4096 0 0 17 50 0 3
352 96
223 96
223 72
0 3 32 0 0 4096 0 0 17 51 0 3
342 109
217 109
217 72
0 4 33 0 0 4096 0 0 17 52 0 3
333 122
211 122
211 72
2 4 30 0 0 8192 0 21 19 0 0 3
310 283
310 347
524 347
0 3 31 0 0 8320 0 0 19 54 0 3
314 248
314 338
524 338
0 2 32 0 0 8320 0 0 19 55 0 3
319 210
319 329
524 329
0 1 33 0 0 8320 0 0 19 56 0 3
326 176
326 320
524 320
0 4 30 0 0 4224 0 0 20 53 0 3
359 283
359 67
528 67
0 3 31 0 0 0 0 0 20 54 0 3
352 248
352 58
528 58
0 2 32 0 0 0 0 0 20 55 0 3
342 210
342 49
528 49
0 1 33 0 0 0 0 0 20 56 0 3
333 176
333 40
528 40
2 4 30 0 0 0 0 21 18 0 0 4
310 283
375 283
375 224
423 224
2 3 31 0 0 0 0 22 18 0 0 4
310 248
380 248
380 215
423 215
2 2 32 0 0 0 0 23 18 0 0 4
309 210
380 210
380 206
423 206
2 1 33 0 0 0 0 24 18 0 0 4
308 176
380 176
380 197
423 197
1 10 34 0 0 8320 0 21 25 0 0 4
274 283
249 283
249 234
236 234
1 11 35 0 0 4224 0 22 25 0 0 4
274 248
244 248
244 225
236 225
1 12 36 0 0 4224 0 23 25 0 0 4
273 210
244 210
244 216
236 216
1 13 37 0 0 8320 0 24 25 0 0 4
272 176
244 176
244 207
236 207
1 2 38 0 0 8320 0 1 25 0 0 4
68 66
142 66
142 198
160 198
1 3 39 0 0 8320 0 2 25 0 0 4
67 114
152 114
152 207
160 207
1 4 40 0 0 4224 0 3 25 0 0 4
68 160
147 160
147 216
160 216
1 5 41 0 0 4224 0 4 25 0 0 4
66 208
152 208
152 225
160 225
1 6 42 0 0 4224 0 5 25 0 0 4
67 257
152 257
152 234
160 234
1 7 43 0 0 4224 0 6 25 0 0 4
65 309
142 309
142 243
160 243
1 8 44 0 0 8320 0 7 25 0 0 4
68 355
147 355
147 252
160 252
1 9 45 0 0 8320 0 8 25 0 0 4
66 402
152 402
152 261
160 261
6
-11 0 0 0 400 0 0 0 0 3 2 1 34
5 Arial
0 0 0 30
875 270 1039 290
882 274 1031 288
30 Decodificador Binario a decima
-11 0 0 0 400 0 0 0 0 3 2 1 34
5 Arial
0 0 0 11
782 266 842 286
786 270 837 284
11 Multiplexor
-11 0 0 0 400 0 0 0 0 3 2 1 34
5 Arial
0 0 0 29
120 139 275 159
127 143 267 157
29 Codificador Decimal a Binario
-11 0 0 0 400 0 0 0 0 3 2 1 34
5 Arial
0 0 0 10
426 137 494 157
430 141 489 155
10 Comparador
-11 0 0 0 400 0 0 0 0 3 2 1 34
5 Arial
0 0 0 7
531 130 589 150
538 134 581 148
7 Sumador
-11 0 0 0 400 0 0 0 0 3 2 1 34
5 Arial
0 0 0 7
527 417 585 437
534 421 577 435
7 Sumador
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
